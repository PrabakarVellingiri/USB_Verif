//===========================================================================
//  CONFIDENTIAL and Copyright (C) 2015 Test and Verification Solutions Ltd
//===========================================================================
//  Contents: 
//   File for class  :   tvs_usb2_ulpi_rx_cmd_test.svh
//
//  Brief description: 
//         This is a test where write_read sequence will execute  
//  Known exceptions to rules:
//    
//============================================================================
//  Author        : 
//  Created on    : 
//  File Id       : 
//============================================================================

`ifndef TVS_USB2_ULPI_RX_CMD_TEST_SVH
`define TVS_USB2_ULPI_RX_CMD_TEST_SVH


///////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////VIRTUAL SEQUENCE//////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
class tvs_usb2_ulpi_rx_cmd_vs#(int DATA_WIDTH =8) extends uvm_sequence#();
 
  ////////////////////////////////////////////////////////////////////////////////
  // Method name         : new 
  // Description         : 
  //                        
  ////////////////////////////////////////////////////////////////////////////////
  function new(string name="tvs_usb2_ulpi_rx_cmd_vs");
    super.new(name);
  endfunction: new
  ////////////////////////////////////////////////////////////////////////////////

  ////////////////////////////////////////////////////////////////////////////////
  //////////////// Register virtual sequence in its virtual sequencer/////////////
  ////////////////////////////////////////////////////////////////////////////////
  `uvm_sequence_utils(tvs_usb2_ulpi_rx_cmd_vs#(DATA_WIDTH),tvs_usb2_virtual_sequencer#(DATA_WIDTH))

  ////////////////////////////////////////////////////////////////////////////////
  ////////////// Respective Sequences needed for the test is included/////////////
  ////////////////////////////////////////////////////////////////////////////////
  // Instance of rx_cmd sequence
  tvs_usb2_host_rx_cmd_sequence#(DATA_WIDTH) rx_cmd_seq;

  ////////////////////////////////////////////////////////////////////////////////
  virtual task pre_body();
    uvm_test_done.raise_objection(this);
  endtask: pre_body
  ////////////////////////////////////////////////////////////////////////////////

  ////////////////////////////////////////////////////////////////////////////////
  // Method name         : Body 
  // Description         : Body of tvs_usb2_ulpi_rx_cmd_seq_vs 
  ////////////////////////////////////////////////////////////////////////////////
  virtual task body();
    begin
      `uvm_do_on_with(rx_cmd_seq,p_sequencer.v_host_sequencer[0],
                     {  linestate_type == IDLE ; 
                        data_type_e    == RX_CMD;    }  )
    end
    #1us;
  endtask: body
                          
 ////////////////////////////////////////////////////////////////////////////////
  virtual task post_body();
    uvm_test_done.drop_objection(this);
  endtask: post_body
  //////////////////////////////////////////////////////////////////////////////// 

endclass : tvs_usb2_ulpi_rx_cmd_vs

///////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////TEST CASE/////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////

class tvs_usb2_ulpi_rx_cmd_test extends tvs_usb2_ulpi_test;

  tvs_usb2_ulpi_rx_cmd_vs#(DATA_WIDTH_SLV) ulpi_rx_cmd_vs;
  ////////////////////////////////////////////////////////////////////////////////
  //////////////////////// Registering the test component/////////////////////////
  //////////////////////////////////////////////////////////////////////////////// 
  `uvm_component_utils(tvs_usb2_ulpi_rx_cmd_test)
  //////////////////////////////////////////////////////////////////////////////// 

  ////////////////////////////////////////////////////////////////////////////////
  // Method name         : new 
  // Description         : Constructor for tvs_usb2_ulpi_rx_cmd_test class. 
  ////////////////////////////////////////////////////////////////////////////////
  function new(string name = "tvs_usb2_ulpi_rx_cmd_test", uvm_component parent=null);
    super.new(name,parent);
  endfunction: new
  ////////////////////////////////////////////////////////////////////////////////
  ////////////////////////////////////////////////////////////////////////////////
  // Method name         : Build 
  // Description         : Configuration of environment as per test case. 
  ////////////////////////////////////////////////////////////////////////////////
  virtual function void build_phase(uvm_phase phase);
    //Create the vip
    super.build_phase(phase);
    // create the object for the sequence 
    ulpi_rx_cmd_vs = tvs_usb2_ulpi_rx_cmd_vs#(.DATA_WIDTH(DATA_WIDTH_SLV))::type_id::create("ulpi_rx_cmd_vs");
  endfunction: build_phase
  ////////////////////////////////////////////////////////////////////////////////
  // Method name         : run_phase 
  // Description         : Start the test sequence
  ///////////////////////////////////////////////////////////////////////////////
  virtual task run_phase(uvm_phase phase);
    uvm_top.print_topology();
    // start the host sequence
    ulpi_rx_cmd_vs.start(usb2_virtual_sequencer);
  endtask: run_phase
  ////////////////////////////////////////////////////////////////////////////////

endclass: tvs_usb2_ulpi_rx_cmd_test

`endif

