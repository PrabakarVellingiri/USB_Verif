package usb_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;

//`include "/tools/questa10_6c/questasim/verilog_src/questa_uvm_pkg-1.2/src/questa_uvm_pkg.sv"
 //import questa_uvm_pkg::*;

`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_declaration.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_seq_item.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_sequences.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_sequencer.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_driver.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_monitor.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_agent.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_arbiter.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_dma.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/scoreboard.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_environment.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_test.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/usb_interface.sv"
`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/USB_VIP/testbench.sv"
//`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/AHB_APB_BRIDGE/TB/test_files/AHB_APB_TEST.sv"
//`include "/Projects/DV_Trainees_Batch2023/devipriya.rajendran/AHB_APB_BRIDGE/TB/AHB_MASTER/AHB_MONITOR.sv"
endpackage

