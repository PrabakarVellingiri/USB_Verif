package usb_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;

`include "usb_declaration.sv"
`include "usb_seq_item.sv"
`include "usb_sequence.sv"
`include "usb_sequencer.sv"
`include "usb_driver.sv"
`include "usb_monitor.sv"
`include "usb_agent.sv"
`include "usb_arbiter.sv"
`include "usb_dma.sv"
`include "usb_scoreboard.sv"
`include "usb_environment.sv"
`include "usb_test.sv"


endpackage

