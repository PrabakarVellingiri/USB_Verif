package WISHBONE_PACKAGE;
`include "uvm_macros.svh"
import uvm_pkg::*;
`include "wb_master_sequence_item.sv"
`include "wb_slave_sequence_item.sv"
`include "wb_master_sequence.sv"
`include "wb_slave_sequence.sv"
`include "wb_master_sequencer.sv"
`include "wb_slave_sequencer.sv"
`include "wb_master_driver.sv"
`include "wb_slave_driver.sv"
`include "wb_master_monitor.sv"
`include "wb_master_agent.sv"
`include "wb_slave_agent.sv"
`include "wb_scoreboard.sv"
`include "wb_environment.sv"
`include "wb_test.sv"

endpackage

