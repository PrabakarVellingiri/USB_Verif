//============================================================================
//  CONFIDENTIAL and Copyright (C) 2015 Test and Verification Solutions Ltd
//============================================================================
//  Contents:
//    File for the list of VIP Files    
//
//  Brief description: 
//    This files contains the list of files in TB Environment included in the
//    compilation/simulation of the design.  
//
//  Known exceptions to rules:
//    
//============================================================================
//  Author        : 
//  Created on    : 
//  File Id       : 
//============================================================================

//----------------------------------------------------------------------------
// UVM Package and Necessary Files 
//----------------------------------------------------------------------------
import uvm_pkg::*;
`include "uvm_macros.svh"
//-----------------------------------------------------------------------------
//--USB2 Package files----------------------------------------------------------
`include "tvs_usb2_top_defines.svh"
import tvs_usb2_device_slave_pkg::*;
import tvs_usb2_host_pkg::*;
import tvs_usb2_env_pkg::*;
import tvs_usb2_test_pkg::*;

//============================================================================
                                                                            
